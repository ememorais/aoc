--Coleção de ROMs que podem ser utilizadas em s1c17_rom.vhd

--ROM Principal
        0  =>  "0000000000000000",  --nop
        1  =>  "1001100100110000",  --ld   %r2, 0x30
        2  =>  "1001101110000111",  --ld   %r7, 0x07
        3  =>  "0000000000000000",  --nop
        4  =>  "0000000000000000",  --nop
        5  =>  "0011100101000111",  --add  %r2, %r7
        6  =>  "1001100000000010",  --ld   %r0, 0x02
        7  =>  "0000000000000000",  --nop
        8  =>  "0011100101010000",  --sub  %r2, %r0
        9 =>  "1001100110000001",   --ld   %r3, 0x01
        10 =>  "0010101100011010",  --ld.a %r6, %r2
        11 =>  "0000000000000000",  --nop
        12 =>  "0000000000000000",  --nop
        13 =>  "0011010101000011",  --cmp.a %r2, %r3
        14 =>  "0000000101001011",  --jpa  %r3

--ROM de teste de ld.a
        0  =>  "0000000000000000",  --nop
        1  =>  "1001100100110000",  --ld   %r2, 0x30
        2  =>  "0000000000000000",  --nop
        3  =>  "0000000000000000",  --nop
        4 =>  "0010101100011010",   --ld.a %r6, %r2

--ROM anterior (lab 5)

        0  =>  "0000000000000000",  --nop
        1  =>  "1001100100110000",  --ld   %r2, 0x30
        2  =>  "1001101110000111",  --ld   %r7, 0x07
        3  =>  "0000000000000000",  --nop
        4  =>  "0000000000000000",  --nop
        5  =>  "0011100101000111",  --add  %r2, %r7
        6  =>  "1001100000000010",  --ld   %r0, 0x02
        7  =>  "0000000000000000",  --nop
        8  =>  "0011100101010000",  --sub  %r2, %r0
        9 =>   "1001100110001000",  --ld   %r3, 0x08
        10 =>  "0010101100011010",  --ld.a %r6, %r2
        11 =>  "0000000000000000",  --nop
        12 =>  "0000000000000000",  --nop
        13 =>  "0011011111000011",  --cmp.a %r7, %r3
        --14 =>  "0011011001000101",  --cmp.a %r4, %r5
        14 =>  "0000000000000000",  --nop
        15 =>  "0000000000000000",  --nop
        16 =>  "0000100001111110",  --jplt -2
        17 =>  "0000000000000000",  --nop
        18 =>  "0000000000000000",  --nop
        19 =>  "0000000101001011",  --jpa  %r3

--Rom lab 6 (conta até 30 e vai somando)

        0  => "0000000000000000", --nop
        1  => "1001100110000000", --ld %r3, 0x00
        2  => "1001101000000000", --ld %r4, 0x00
        3  => "1001101010000001", --ld %r5, 0x01
        4  => "1001101100011110", --ld %r6, 0x30
        5  => "0011101001000011", --add %r4, %r3
        6  => "0011100111000101", --add %r3, %r5 (r3 + 1)
        7  => "0000000000000000", --nop
        8  => "0000000000000000", --nop
        9  => "0011010111000110", --cmp %r3, %r6 (r3, 30)
        10 => "0000000000000000", --nop
        11 => "0000000000000000", --nop
        12 => "0000100001110111", --jplt -9
        13 => "0000000000000000", --nop
        14 => "0000000000000000", --nop
        15 => "0010101010011100", --ld %r5, r4