

        --FIM DO FOR